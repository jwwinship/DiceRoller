module d_bounce(



);


endmodule