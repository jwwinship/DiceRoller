module RNG(input  wire clk,
              input  wire reset,
              input  wire start,
              output wire [31:0] result,
	      output wire done);
   
   
   
endmodule
